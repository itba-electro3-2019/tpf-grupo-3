localparam LEFT_START = 10'd50;
localparam RIGHT_START = 10'd590;
localparam TOP = 10'd20;
localparam BOT = 10'd25;
localparam W = 10'd5;
localparam SPACE = 10'd5;