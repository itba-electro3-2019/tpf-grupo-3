localparam X_GMV_LEFT1 = 0;
localparam X_GMV_LEFT2 = 320;
localparam X_GMV_RIGHT1 = 320;
localparam X_GMV_RIGHT2 = 640;
localparam Y_GMV_TOP = 0;
localparam Y_GMV_BOT = 480;
localparam Y_FLOOR = 475;
localparam Y_CEIL = 5;
localparam X_LWALL = 5;
localparam X_RWALL = 635;
localparam BALL_H = 10;
localparam BALL_W = 10;
localparam PAD_H = 100;
localparam ALT_PAD_H = 150;
localparam ALT2_PAD_H = 60;
localparam PAD_W = 12;
localparam Y_BALL_VEL = 2;
localparam X_BALL_VEL = 2;
localparam ALT_X_BALL_VEL = 3;
localparam Y_PAD_VEL = 2;
localparam ALT_Y_PAD_VEL = 4;
localparam X_PAD_VEL = 2;
localparam X_BALL_DEF = 315;
localparam Y_BALL_DEF = 235;
localparam X_PADA_DEF = 20;
localparam X_PADB_DEF = 610;
localparam Y_PAD_DEF = 200;
localparam BALL_DIR_DEF = 1;
localparam DEF_SCR = 0;
localparam LEFT = 0;
localparam UP = 0;
localparam DOWN = 1;
localparam RIGHT = 1;
localparam NORMAL = 0;
localparam LONG_PAD = 1;
localparam QUICK_PAD = 2;
localparam QUICK_BALL = 3;
localparam SMALL_PAD = 4;
localparam INVERTED_PAD = 5;
localparam FLICK_PAD = 6;
localparam POWER_UP_H = 17;
localparam POWER_UP_W = 17;
localparam PADBUZZ = 3;
localparam WALLBUZZ = 6;
localparam POWER_OFF_COUNT = 1300;
localparam POWER_SPAWN_COUNT = 2000;