module PaddleCollisionController(

);




endmodule